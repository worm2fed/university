module segmentdisplay (x1, x2, x3, x4, a, b, c, d, e, f, g);
	input x1, x2, x3, x4;
	output a, b, c, d, e, f, g;
	
	// x1 x2 x3 x4 | a b c d e f g			 	a		    b			c		    d			e		    f			g
	// ------------|--------------			-----------------   -----------------   -----------------   -----------------   -----------------   -----------------   -----------------
	// 0  0  0  0  | 1 1 1 1 1 1 0			| + |   | + | + |   | + | + |   | + |   | + | + |   | + |   | + |   | + | + |   | + |   | + | + |   | + | + | + | + |   |   | + |   | + |   
	// 0  0  0  1  | 0 1 1 0 0 0 0			-----------------   -----------------   -----------------   -----------------   -----------------   -----------------   -----------------
	// 0  0  1  0  | 1 1 0 1 1 0 1			|   | + |   | + |   | + |   | + | + |   | + | + | + | + |   |   | + | + |   |   |   |   | + |   |   |   | + |   | + |   |   | + | + | + |   
	// 0  0  1  1  | 1 1 1 1 0 0 1			-----------------   -----------------   -----------------   -----------------   -----------------   -----------------   -----------------
	// 0  1  0  0  | 0 1 1 0 0 1 1			| + | + | + |   |   | + | + |   |   |   | + | + |   | + |   | + |   |   | + |   |   |   | + | + |   |   |   | + | + |   | + |   | + | + |   
	// 0  1  0  1  | 1 0 1 1 0 1 1			-----------------   -----------------   -----------------   -----------------   -----------------   -----------------   -----------------
	// 0  1  1  0  | 1 0 1 1 1 1 1			| + | + | + | + |   | + |   |   | + |   |   | + |   | + |   | + | + | + |   |   | + | + | + | + |   |   | + | + | + |   | + | + | + | + |   
	// 0  1  1  1  | 1 1 1 0 0 0 0			-----------------   -----------------   -----------------   -----------------   -----------------   -----------------   -----------------
	// 1  0  0  0  | 1 1 1 1 1 1 1			
	// 1  0  0  1  | 1 1 1 0 0 1 1			a = x3!x4 + x1x2x3 + !x1x3x4 + !x1x2x4 + !x2!x3!x4 + x1!x3!x4 + x1!x2!x3
	// 1  0  1  0  | 1 1 1 0 1 1 1			b = !x1!x3!x4 + x1!x3x4 + x1!x2!x4 + !x1x3x4 + !x1!x2
	// 1  0  1  1  | 0 0 1 1 1 1 1			c = !x1x3x4 + !x3x4 + !x2!x3 + !x1x2 + x1!x2
	// 1  1  0  0  | 1 0 0 1 1 1 0			d = !x1!x2!x4 + !x2x3x4 + x2x3!x4 + x2!x3x4 + x1x2!x3 + !x2!x3!x4
	// 1  1  0  1  | 0 1 1 1 1 0 1			e = !x2!x4 + x1x2 + x1x3 + x3!x4
	// 1  1  1  0  | 1 0 0 1 1 1 1			f = !x1x2!x3 + x2x3!x4 + x1x3 + !x3!x4 + x1!x2
	// 1  1  1  1  | 1 0 0 0 1 1 1			g = !x1x2!x3 + x1!x2!x3 + x1x4 + x3!x4 + !x1!x2x3
	
	assign a = x3 & !x4 | x1 & x2 & x3 | !x1 & x3 & x4 | !x1 & x2 & x4 | !x2 & !x3 & !x4 | x1 & !x3 & !x4 | x1 & !x2 & !x3;
	assign b = !x1 & !x3 & !x4 | x1 & !x3 & x4 | x1 & !x2 & !x4 | !x1 & x3 & x4 | !x1 & !x2;
	assign c = !x1 & x3 & x4 | !x3 & x4 | !x2 & !x3 | !x1 & x2 | x1 & !x2;
	assign d = !x1 & !x2 & !x4 | !x2 & x3 & x4 | x2 & x3 & !x4 | x2 & !x3 & x4 | x1 & x2 & !x3 | !x2 & !x3 & !x4;
	assign e = !x2 & !x4 | x1 & x2 | x1 & x3 | x3 & !x4;
	assign f = !x1 & x2 & !x3 | x2 & x3 & !x4 | x1 & x3 | !x3 & !x4 | x1 & !x2;
	assign g = !x1 & x2 & !x3 | x1 & !x2 & !x3 | x1 & x4 | x3 & !x4 | !x1 & !x2 & x3;
endmodule

